module top_module(input in, output out);
	assign out = in; // creates a wire from input to output
endmodule